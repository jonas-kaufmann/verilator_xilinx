`ifdef verilator3
`else
`timescale 1 ps / 1 ps
`endif
//
// RAM512X1S primitive for Xilinx FPGAs
// Compatible with Verilator tool (www.veripool.org)
// Copyright (c) 2019-2022 Frédéric REQUIN
// License : BSD
//

/* verilator coverage_off */
/* verilator tracing_off */
module RAM512X1S
#(
    parameter [511:0] INIT = 512'h0,
    parameter   [0:0] IS_WCLK_INVERTED = 1'b0
)
/* verilator tracing_on */
(
    // Write clock
    input  wire       WCLK,
    // Write enable
    input  wire       WE,
    // Read / Write address
    input  wire [8:0] A,
    // Data in
    input  wire       D,
    // Data out
    output wire       O
);
/* verilator tracing_off */
    // 512 x 1-bit Select RAM
    reg  [511:0] _r_mem;
    
    // Power-up value
    initial begin : INIT_STATE
        _r_mem = INIT;
    end
    
    // Synchronous memory write
    generate
        if (IS_WCLK_INVERTED) begin : GEN_WCLK_NEG
            always @(negedge WCLK) begin : MEM_WRITE
            
                if (WE) begin
                    _r_mem[A] <= D;
                end
            end
        end
        else begin : GEN_WCLK_POS
            always @(posedge WCLK) begin : MEM_WRITE
            
                if (WE) begin
                    _r_mem[A] <= D;
                end
            end
        end
    endgenerate
    
    // Asynchronous memory read
    assign O = _r_mem[A];

endmodule
/* verilator coverage_on */
